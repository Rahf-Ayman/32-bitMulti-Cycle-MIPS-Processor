library ieee;
use ieee.std_logic_1164.all;

entity connection is
	port (
	CLK : in std_logic;
	reset : in std_logic
	);
end connection;

architecture behavior of connection is
-- component of register
	-- here
--

-- component of dataflow
	-- here
--

-- component of control unit
	-- here
--

-- internal signal
	-- here
--
begin
-- port map of register
	-- here
--

-- port map of dataflow
	-- here
--

-- port map of control unit
	-- here
--	
end behavior;
	